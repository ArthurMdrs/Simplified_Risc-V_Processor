module data_mem_vc #(
    int AWIDTH = 3,
    int DWIDTH = 8
) (
    input  logic [DWIDTH-1:0] rdata,
    input  logic [DWIDTH-1:0] wdata,
    input  logic [AWIDTH-1:0] addr,
    input  logic              wen,
    input  logic              clk,
    input  logic              rst_n
);    

`ifdef SVA_ON

// Defaults
default clocking def_clk @(posedge clk); 
endclocking

default disable iff (!rst_n);

// Aux code
bit write_happened;
always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n)
        write_happened <= 0;
    else if (wen)
        write_happened <= 1;
end



// Properties
property SIGNAL_CAN_BE_VALUE (signal, value);
    (signal == value);
endproperty

property NO_RDATA_WO_WRITE (rdata);
    (rdata != 0) |-> (write_happened);
endproperty



// Assertions
AST_NO_RDATA_WO_WRITE: assert property (NO_RDATA_WO_WRITE(rdata));



// Covers
generate
    for (genvar i = 0; i < DWIDTH; i++) begin
        COV_RDATA_CAN_BE_VAL: cover property (SIGNAL_CAN_BE_VALUE(rdata, 2**i-1));
    end
endgenerate



`ifndef SIM

// Data integrity check (NDC only possible in formal!)

bit [AWIDTH-1:0] addr_ndc; // Non-deterministic constant
bit [DWIDTH-1:0] xptd_data; // Expected data
bit wr_to_addr_ndc; // Write to addr_ndc location
always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        xptd_data <= '0;
        wr_to_addr_ndc <= 0;
    end else if (wen && addr == addr_ndc) begin
        xptd_data <= wdata;
        wr_to_addr_ndc <= 1;
    end
end

property DATA_INTEGRITY (raddr, rdata);
    (wr_to_addr_ndc && raddr == addr_ndc) |-> (rdata == xptd_data);
endproperty 

AST_DATA_INTEGRITY1: assert property (DATA_INTEGRITY(addr, rdata));

ASM_ADDR_NDC_NOT_0: assume property (addr_ndc != '0);
ASM_ADDR_NDC_CONST: assume property (addr_ndc == $past(addr_ndc));

`endif
    
`endif

endmodule